`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/21/2022 01:20:59 AM
// Design Name: 
// Module Name: test_env
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_env(
    input clk,
    input [4:0] btn,
    input [15:0] sw,
    output [15:0] led,
    output [3:0] an,
    output [6:0] cat
    );
endmodule
